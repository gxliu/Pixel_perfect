`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:03:02 11/08/2012 
// Design Name: 
// Module Name:    dcm_cust_clk 
//////////////////////////////////////////////////////////////////////////////////
module dcm_cust_clk(
    );


endmodule
